library ieee;
use ieee.std_logic_1164.all;

entity practica_1 is
port (x: in std_logic_vector(3 downto 0);
 z: out std_logic_vector(1 downto 0));
end practica_1;


architecture estructural_deco of practica_1 is
signal a: std_logic_vector(2 downto 0);
signal b: std_logic_vector(7 downto 0);

begin 

a(0) <= x (1);
a(1) <= x (2);
a(2) <= x (3);

deco: entity work.deco3a8(funcional) port map ('1',a,b);
z(0) <= (b(1) or (b(2) and x(0)) or (b(3) and x(0)) or (b(5) and x(0)) or (b(6) and x(0)));
z(1) <= (b(0) or b(1) or (b(2) and x(0)) or (b(4) and (not x(0))) or (b(6) and x(0)));
end estructural_deco;
